LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
PACKAGE seven_segment_display_package IS
COMPONENT seven_segment_display
PORT ( W,X ,Y,Z       : IN STD_LOGIC;
      A,B,C,D,E,F,G   : OUT STD_LOGIC);
END COMPONENT ;
END seven_segment_display_package ;
