Library ieee;
USE ieee.std_logic_1164.all;
ENTITY seven_segment_display IS
PORT (W,X,Y,Z         : IN STD_LOGIC;
      A,B,C,D,E,F,G   : OUT STD_LOGIC);
END seven_segment_display;
ARCHITECTURE LogicFunc OF seven_segment_display IS
BEGIN
A <= (X AND NOT Y AND NOT Z) OR (W AND X AND NOT Y) OR (NOT W AND NOT X AND NOT Y AND Z) OR (W AND NOT X AND Y AND Z);
B <= (X AND Y AND NOT Z) OR (W AND X AND Y) OR (W AND Y AND Z) OR (W AND X AND NOT Z) OR (NOT W AND X AND NOT Y AND Z);
C <= (NOT W AND NOT X AND Y AND NOT Z) OR (W AND X AND NOT Z) OR (W AND X AND Y);
D <= (NOT X AND NOT Y AND Z) OR (NOT W AND X AND NOT Y AND NOT Z) OR (X AND Y AND Z) OR (W AND NOT X AND Y AND NOT Z);
E <= (NOT W AND Z) OR (NOT W AND X AND NOT Y) OR (NOT X AND NOT Y AND Z);
F <= (NOT W AND NOT X AND Z) OR (NOT W AND NOT X AND Y) OR (NOT W AND Y AND Z) OR (W AND X AND NOT Y);
G <= (NOT W AND NOT X AND NOT Y) OR (NOT W AND X AND Y AND Z);
END LogicFunc;
