Library ieee;
USE ieee.std_logic_1164.all;
ENTITY GOAL_two IS
PORT (W,X,Y,Z,w1,x1,y1,z1         : IN STD_LOGIC;
      A,B,C,D,E,F,G,a1,b1,c1,d1,e1,f1,g1   : OUT STD_LOGIC);
END GOAL_two;
ARCHITECTURE LogicFunc OF GOAL_twos IS
BEGIN
A <= (X AND NOT Y AND NOT Z) OR (W AND X AND NOT Y) OR (NOT W AND NOT X AND NOT Y AND Z) OR (W AND NOT X AND Y AND Z);
B <= (X AND Y AND NOT Z) OR (W AND X AND Y) OR (W AND Y AND Z) OR (W AND X AND NOT Z) OR (NOT W AND X AND NOT Y AND Z);
C <= (NOT W AND NOT X AND Y AND NOT Z) OR (W AND X AND NOT Z) OR (W AND X AND Y);
D <= (NOT X AND NOT Y AND Z) OR (NOT W AND X AND NOT Y AND NOT Z) OR (X AND Y AND Z) OR (W AND NOT X AND Y AND NOT Z);
E <= (NOT W AND Z) OR (NOT W AND X AND NOT Y) OR (NOT X AND NOT Y AND Z);
F <= (NOT W AND NOT X AND Z) OR (NOT W AND NOT X AND Y) OR (NOT W AND Y AND Z) OR (W AND X AND NOT Y);
G <= (NOT W AND NOT X AND NOT Y) OR (NOT W AND X AND Y AND Z);

a1 <= (x1 AND NOT y1 AND NOT z1) OR (w1 AND x1 AND NOT y1) OR (NOT w1 AND NOT x1 AND NOT y1 AND z1) OR (w1 AND NOT x1 AND y1 AND z1);
b1 <= (x1 AND y1 AND NOT z1) OR (w1 AND x1 AND y1) OR (w1 AND y1 AND z1) OR (w1 AND x1 AND NOT z1) OR (NOT w1 AND x1 AND NOT y1 AND z1);
c1 <= (NOT w1 AND NOT x1 AND y1 AND NOT z1) OR (w1 AND x1 AND NOT z1) OR (w1 AND x1 AND y1);
d1 <= (NOT x1 AND NOT y1 AND z1) OR (NOT w1 AND x1 AND NOT y1 AND NOT z1) OR (x1 AND y1 AND z1) OR (w1 AND NOT x1 AND y1 AND NOT z1);
e1 <= (NOT w1 AND z1) OR (NOT w1 AND x1 AND NOT y1) OR (NOT x1 AND NOT y1 AND z1);
f1 <= (NOT w1 AND NOT x1 AND z1) OR (NOT w1 AND NOT x1 AND y1) OR (NOT w1 AND y1 AND z1) OR (w1 AND x1 AND NOT y1);
g1 <= (NOT w1 AND NOT x1 AND NOT y1) OR (NOT w1 AND x1 AND y1 AND z1);
END LogicFunc;