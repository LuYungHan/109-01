LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
PACKAGE fulladd_package IS
COMPONENT fulladd
PORT ( Cin, x, y : IN STD_LOGIC ;
s, Cout : OUT STD_LOGIC ) ;
END COMPONENT ;
END fulladd_package ;
